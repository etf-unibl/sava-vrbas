-----------------------------------------------------------------------------
-- Faculty of Electrical Engineering
-- PDS 2022
-- https://github.com/knezicm/sava-vrbas/
-----------------------------------------------------------------------------
--
-- unit name:    24-BIT BUFFER VUNIT TESTBENCH
--
-- description:
--
--  This file implements 24-bit buffer testbench, following  VUnit testbench form.
--
-----------------------------------------------------------------------------
-- Copyright (c) 2022 Faculty of Electrical Engineering
-----------------------------------------------------------------------------
-- The MIT License
-----------------------------------------------------------------------------
-- Copyright 2022 Faculty of Electrical Engineering
--
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the "Software"),
-- to deal in the Software without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Software, and to permit persons to whom
-- the Software is furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
-- THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE
-----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_1164;
use ieee.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_context;

use vunit_lib.run_pkg.all;
use vunit_lib.check_pkg.all;

library common_lib;

entity tb_example is
  generic (runner_cfg : string);
end entity;

architecture tb of tb_example is
  signal write_enable_i : std_logic;
  signal data_i : std_logic_vector(23 downto 0);
  signal data_o : std_logic_vector(23 downto 0) := (others => '0');

begin
  invdut : entity common_lib.buffer24
    port map(
      write_enable_i => write_enable_i,
      data_i => data_i,
      data_o => data_o);

  clock_stimulus : process
  begin
    write_enable_i <= '1';
    wait for 100 ns;
    write_enable_i <= '0';
    wait for 100 ns;
  end process;

  test_runner : process
  begin
    test_runner_setup(runner, runner_cfg);

    while test_suite loop

      if run("check_input_no_enable") then
        info("Performing first test");
        data_i <= std_logic_vector'("011001101000110010011010");
        wait for 1000 ns;
        write_enable_i <= '0';
        -- This test passes
        check_equal(data_o, std_logic_vector'("000000000000000000000000"));

      elsif run("check_input_with_enable") then
        info("Performing second test");
        write_enable_i <= '1';
        data_i <= std_logic_vector'("011001101000110010011010");
        wait for 1000 ns;
        -- This test constantly fails, output is unable to change its value to data_i
        check_equal(data_o, std_logic_vector'("011001101000110010011010"));
      end if;
      test_runner_cleanup(runner);
    end loop;

  end process;
end architecture;